module logic_gates( input logic and,)