library verilog;
use verilog.vl_types.all;
entity triggers_tb is
end triggers_tb;
