`timescale 1 ns/10ps // time-unit = 1ns, precision = 10 ps

module silyfunction_tb();
    reg a, b, c;
    wire y;

    sillyfunction dut (.a(a), .b(b), .c(c), .y(y));

    initial begin
      a = 0; b = 0; c = 0; #10;
      c = 1; #10
      b = 1; c =0; #10;
      c = 1; #10 
      a = 1; b = 0; c = 0; #10;
    end
endmodule